module iinv(output z, input a);
	assign z = ~a;
endmodule 
