module example(/*AUTOARG*/);
	input i;
	output o;
/*AUTOINPUT*/
/*AUTOOUTPUT*/
/*AUTOREG*/
inst inst (/*AUTOINST*/);
always@(/*AUTOSENSE*/) begin
o = i;
end
endmodule
