module bbuf(output z, input a);
	assign z = a;
endmodule 
