module aand(output z, input a, input b);
	assign z = a & b;
endmodule
