module inst(
	input lower_ina,
	input lower_inb,
	output lower_out
);

endmodule
